//transcation for and gate

class and_transaction;
	rand bit a_i, b_i;
	bit y_o;
endclass


