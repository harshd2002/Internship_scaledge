class ram_base_test;

  //take handle of verification environment class
  
  //declare all interface 
  
   //take new method (only for virtual interface)
   
   //call environment method here as needed
   task build_and_run();
    :
endtask
     
  
endclass