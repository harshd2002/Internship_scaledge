////////////////////////////////////////////////////////////////////////////////////////////////////
//
//
//Header
//
//
////////////////////////////////////////////////////////////////////////////////////////////////////

//APB global variables declaration

`ifndef APB_DEFINE
`define APB_DEFINE

`define DRV_PATH  vintf.apb_mp_drv.apb_cb_drv
`define MON_PATH  vintf.apb_mp_mon.apb_cb_mon

`endif
