//No we cannot access local property of parent class directly in child class

