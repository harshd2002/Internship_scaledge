//randomize array of size 5 to 10 having values in ascending and descending order

class order_arr;
	rand byte arr_a[];
	rand byte arr_d[];
endclass

module que_8();

endmodule
