////////////////////////////////////////////////////////////////////////////////////////////////////
//
//
//Header
//
//
////////////////////////////////////////////////////////////////////////////////////////////////////

//APB generator class

`define DRV_PATH vintf.apb_mp_drv.apb_cb_drv
`define MON_PATH vintf.apb_mp_mon.apb_cb_mon

//enum type variable to select operation type
typedef enum {PWRITE, PREAD} operation;
