class ram_env;

  //take handles of all verification sub component
  
  //declare all mailboxs
  
  //declare all interface 
  
   //take new method (only for virtual interface)
   
   //create all the component in this method
   task build();
     :
  endtask
  
  //call all sub verif component run task in parallel
  task run();
  :
  endtask
  
endclass
   
  