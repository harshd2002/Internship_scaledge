module decoder_5x32(input wire enbl,
	input wire [4:0] inp,
	output wire [31:0] out
	);
	
	reg [31:0] out_r;

	always @(*) begin

		if(enbl) begin

			case(

		end

	end

endmodule
