//RAM files are included

package pkg_files;
	event item_done;
	`include "ram_trans.sv"
	`include "ram_gen.sv"
	`include "ram_drv.sv"
	`include "ram_mon.sv"
	`include "ram_pred.sv"
	`include "ram_scrbd.sv"
	`include "ram_env.sv"
	`include "ram_test.sv"
endpackage
