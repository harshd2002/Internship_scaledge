//generate prime number

class prime_class;
	
endclass
