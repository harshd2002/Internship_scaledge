package pkg_files;

  `include "global_define.sv"
  `include "transaction.sv"
  `include "generator.sv"
  `include "gen_sanity.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "predictor.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "test.sv"

endpackage
