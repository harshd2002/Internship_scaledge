

`include "ram_interface.sv"
package ram_pkg;
 event item_done_ev;
  //`include "ram_defines.sv
  //`include "ram_trans.sv
  //add all file till test, don't miss the order
  
endpackage