

module ram_tb_top();

  //generate clock
  
  //take instance of actual interface
  
  
  //take intance of test class
  
  
  //instantiate design
  ram DUT (.clk(clk),
           .rst(inf.rst),
		   .wr_enb(inf.we)
  
  //
  initial
    //create test
	//call require test method
	
	:

endmodule