package pkg_files;

  `include "global_define.sv"
  `include "transaction.sv"
  `include "generator.sv"
  `include "gen_sanity.sv"
  `include "gen_sel_0.sv"
  `include "gen_sel_1.sv"
  `include "gen_sel_2.sv"
  `include "gen_sel_3.sv"
  `include "gen_sel_4.sv"
  `include "gen_sel_5.sv"
  `include "gen_sel_6.sv"
  `include "gen_inbet_reset.sv"
  `include "gen_invalid_sel.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "predictor.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "test.sv"

endpackage
