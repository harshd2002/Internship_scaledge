//randomize a variable
//values should be greator than 50
//override the constraint and store values less than 50

class question22b;
	rand int a;
	constraint c1 {
		a > 50;
	}

endclass

module constraint_override();

endmodule
