// AND gate monitor class

class and_mon;

endclass
