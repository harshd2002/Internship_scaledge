class ram_scoreboard;

  //take transation handles
  
  //declare mailbox
  
  //take new method
  
  
  task run();
   repeat(10) begin
    //collect data from all mailbox
	//compare act and exp and log the results
   end
  endtask
    
  //description
 task check_data(ram_trans act_trans, ram_trans exp_trans);
  
 endtask
  
 endclass